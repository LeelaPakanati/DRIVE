//COM Stage*******************************************************
reorderbuf rob(
	.clk(clk),
	.reset(reset),
	.dp1(~stall_DP & ~kill_DP & ~inv1_id),
	.dp1_addr(dst1_renamed),
	.pc_dp1(pc_id),
	.storebit_dp1(inst1_id[6:0] == `RV32_STORE ? 1'b1 : 1'b0),
	.dstvalid_dp1(wr_reg_1_id),
	.dst_dp1(rd_1_id),
	.bhr_dp1(bhr_id),
	.isbranch_dp1(req1_branch),
	.dp2(~stall_DP & ~kill_DP & ~inv2_id),
	.dp2_addr(dst2_renamed),
	.pc_dp2(pc_id + 4),
	.storebit_dp2(inst2_id[6:0] == `RV32_STORE ? 1'b1 : 1'b0),
	.dstvalid_dp2(wr_reg_2_id),
	.dst_dp2(rd_2_id),
	.bhr_dp2(bhr_id),
	.isbranch_dp2(req2_branch),
	.exfin_alu1(robwe_alu1),
	.exfin_alu1_addr(buf_rrftag_alu1),
	.exfin_alu2(robwe_alu2),
	.exfin_alu2_addr(buf_rrftag_alu2),
	.exfin_mul(robwe_mul),
	.exfin_mul_addr(buf_rrftag_mul),
	.exfin_ldst(robwe_ldst),
	.exfin_ldst_addr(wrrftag_ldst),
	.exfin_branch(robwe_branch),
	.exfin_branch_addr(buf_rrftag_branch),
	.exfin_branch_brcond(brcond),
	.exfin_branch_jmpaddr(jmpaddr_taken),
	.exfin_C1(robwe_C1),
	.exfin_C1_addr(buf_rrftag_C1),
	.exfin_C2(robwe_C2),
	.exfin_C2_addr(buf_rrftag_C2),

	.comptr(comptr),
	.comptr2(comptr2),
	.comnum(comnum),
	.stcommit(stcommit),
	.arfwe1(arfwe1),
	.arfwe2(arfwe2),
	.dstarf1(dstarf1),
	.dstarf2(dstarf2),
	.pc_combranch(pc_combranch),
	.bhr_combranch(bhr_combranch),
	.brcond_combranch(brcond_combranch),
	.jmpaddr_combranch(jmpaddr_combranch),
	.combranch(combranch),
	.dispatchptr(rrfptr),
	.rrf_freenum(freenum),
	.prmiss(prmiss)
	);