rs_requestgenerator rs_reqgen(
	.rsent_1(rs_ent_1_id),
	.rsent_2(rs_ent_2_id),
	.req1_alu(req1_alu),
	.req2_alu(req2_alu),
	.req_alunum(req_alunum),
	.req1_branch(req1_branch),
	.req2_branch(req2_branch),
	.req_branchnum(req_branchnum),
	.req1_mul(req1_mul),
	.req2_mul(req2_mul),
	.req_mulnum(req_mulnum),
	.req1_ldst(req1_ldst),
	.req2_ldst(req2_ldst),
	.req_ldstnum(req_ldstnum),
	.req1_C1(req1_C1),
	.req2_C1(req2_C1),
	.req_C1num(req_C1num),
	.req1_C2(req1_C2),
	.req2_C2(req2_C2),
	.req_C2num(req_C2num)
	);