`define	RS_ENT_C1 5
`define	RS_ENT_C2 6


`define C1_ENT_SEL 1
`define C1_ENT_NUM 2
`define C2_ENT_SEL 1
`define C2_ENT_NUM 2

`define C1	0
`define C2	1